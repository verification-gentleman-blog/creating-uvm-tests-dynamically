module top;

  import uvm_pkg::*;


  initial
    run_test("test_that_executes_some_sequence");

endmodule
