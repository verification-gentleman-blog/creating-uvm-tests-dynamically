module top;

  import uvm_pkg::*;


  initial
    run_test();

endmodule
