class wrapper_for_test_that_executes_some_sequence_using_param
    extends uvm_component_registry #(test_that_executes_sequence_via_param #(some_sequence), "test_that_executes_some_sequence_using_param");
endclass
