package generic_test_builder;

  import uvm_pkg::*;
  `include "uvm_macros.svh"


  `include "test_that_executes_sequence.svh"
  `include "wrapper_for_test_that_executes_sequence.svh"
  `include "test_builder.svh"

endpackage
